module keyboard
